module VGA_overlay (
    input               iCLK,
    input               iRST_N,
    input               iVideo_On,

    input       [10:0]  iVga_x,
    input       [10:0]  iVga_y,

    input       [9:0]   iRed,
    input       [9:0]   iGreen,
    input       [9:0]   iBlue,

    output reg  [9:0]   oRed,
    output reg  [9:0]   oGreen,
    output reg  [9:0]   oBlue
);

	// VIDEO REGION
	parameter WIDTH 	 = 600;
	parameter HEIGHT   = 430;
	parameter VIDEO_X0 = (640 - WIDTH) / 2;
	parameter VIDEO_Y0 = 120;	// 20 px below text
	
	wire video_region  = (iVga_x >= VIDEO_X0 & iVga_x < (VIDEO_X0 + WIDTH) &
								 iVga_y >= VIDEO_Y0 & iVga_y < (VIDEO_Y0 + HEIGHT));
								 
    // ----------------------
    // Parameters
    // New character size: 16x32 (2x scaled from 8x16)
    // ----------------------
    parameter WHITE = 10'h3FF;
    parameter BLACK = 10'h000;
	 parameter RED   = 10'hF00;
	 parameter GREEN = 10'h0F0;
	 
	 
    parameter CHAR_WIDTH = 16;  // Doubled from 8
    parameter CHAR_HEIGHT = 32; // Doubled from 16
	 
	 parameter CHAR_WIDTH2 = 32;  // Doubled from 8
    parameter CHAR_HEIGHT2 = 64; // Doubled from 16

    // Text strings
    localparam VIDEO_ON_TEXT = "INTRUDER";
    localparam VIDEO_OFF_TEXT = "ARMED";

    localparam VIDEO_ON_LEN  = 8;
    localparam VIDEO_OFF_LEN = 5;

    // ----------------------
    // Compute text position (centered - uses new CHAR_WIDTH and CHAR_HEIGHT)
    // ----------------------
    wire [10:0] TEXT_X0  = (640 - (VIDEO_ON_LEN * CHAR_WIDTH)) / 2;
    wire [10:0] TEXT_Y0  = 50;

    wire [10:0] TEXT_X02 = (640 - (VIDEO_OFF_LEN * CHAR_WIDTH2)) / 2;
    wire [10:0] TEXT_Y02 = (480 - (CHAR_HEIGHT2)) / 2;

    // ----------------------
    // Determine if pixel is in text region
    // ----------------------
    wire in_text_on  = (iVga_x >= TEXT_X0  && iVga_x <  TEXT_X0 + VIDEO_ON_LEN  * CHAR_WIDTH) &&
                       (iVga_y >= TEXT_Y0  && iVga_y < TEXT_Y0  + CHAR_HEIGHT);

    wire in_text_off = (iVga_x >= TEXT_X02 && iVga_x < TEXT_X02 + VIDEO_OFF_LEN * CHAR_WIDTH2) &&
                       (iVga_y >= TEXT_Y02 && iVga_y < TEXT_Y02 + CHAR_HEIGHT2);

    // ----------------------
    // Compute character index & pixel inside character (uses new 16x32 bounds)
    // ----------------------
    // char_x_full (0 to 15)
    wire [3:0] char_x_full = (iVga_x - TEXT_X0)  % CHAR_WIDTH;
    // char_y_full (0 to 31)
    wire [4:0] char_y_full = (iVga_y - TEXT_Y0)  % CHAR_HEIGHT;

    // Low-resolution 8x16 coordinates for ROM lookup (Pixel Doubling)
    // By using bits [3:1] of char_x_full, the LSB (bit 0) is ignored, doubling the width.
    wire [2:0] char_x_low = char_x_full[3:1]; // 8-pixel index (0 to 7)
    // By using bits [4:1] of char_y_full, the LSB (bit 0) is ignored, doubling the height.
    wire [3:0] char_y_low = char_y_full[4:1]; // 16-row index (0 to 15)

	 
    // Character index is based on the 16-pixel width
    wire [2:0] char_idx = (iVga_x - TEXT_X0) / CHAR_WIDTH;
	 
	 
	 
	 
	 
	 
	 wire [4:0] char_x_full2 = (iVga_x - TEXT_X02)  % CHAR_WIDTH2;
    // char_y_full (0 to 31)
    wire [5:0] char_y_full2 = (iVga_y - TEXT_Y02) % CHAR_HEIGHT2;

    // Low-resolution 8x16 coordinates for ROM lookup (Pixel Doubling)
    // By using bits [3:1] of char_x_full, the LSB (bit 0) is ignored, doubling the width.
    wire [2:0] char_x_low2 = char_x_full2[4:2]; // 8-pixel index (0 to 7)
    // By using bits [4:1] of char_y_full, the LSB (bit 0) is ignored, doubling the height.
    wire [3:0] char_y_low2 = char_y_full2[5:2]; // 16-row index (0 to 15)

    // Character index is based on the 16-pixel width
    wire [2:0] char_idx2 = (iVga_x - TEXT_X02) / CHAR_WIDTH2;

	 
	 
	 
    // ----------------------
    // Select ASCII code for current character (same logic)
    // ----------------------
    reg [6:0] ascii_code;
	 reg [6:0] ascii_code2;
	 
    always @* begin
		ascii_code = 7'h20;
		ascii_code2 = 7'h20;
		
        if(iVideo_On && in_text_on) begin
            case(char_idx)
                0: ascii_code = "I";
                1: ascii_code = "N";
                2: ascii_code = "T";
                3: ascii_code = "R";
                4: ascii_code = "U";
                5: ascii_code = "D";
                6: ascii_code = "E";
                7: ascii_code = "R";
                default: ascii_code = 7'h20;
            endcase
        end
        else if(!iVideo_On && in_text_off) begin
            case(char_idx2)
                0: ascii_code2 = "A";
                1: ascii_code2 = "R";
                2: ascii_code2 = "M";
                3: ascii_code2 = "E";
                4: ascii_code2 = "D";
                default: ascii_code2 = 7'h20;
            endcase
        end
    end

    // ----------------------
    // ASCII ROM address and output
    // Use the low-resolution row for addressing
    // ----------------------
    wire [10:0] rom_addr = {ascii_code, char_y_low};
	 wire [10:0] rom_addr2 = {ascii_code2, char_y_low2}; 
    wire [7:0] rom_out;
	 wire [7:0] rom_out2;
	 
    ascii_rom (
        .addr(rom_addr),
        .data(rom_out)
    );
	 
	 ascii_rom (
        .addr(rom_addr2),
        .data(rom_out2)
    );
	 
	 

    // rom_out[7 - char_x_low] gets the pixel state for the low-res 8x16 character.
    // This state is then used across 2x2 screen pixels.
    wire pixel_on = iVideo_On && in_text_on && rom_out[7 - char_x_low];
	 
											
	 wire pixel_on2 = !iVideo_On && in_text_off && rom_out2[7 - char_x_low2];

    // ----------------------
    // VGA output (remains the same)
    // ----------------------
    always @(posedge iCLK) begin
        if (!iRST_N) begin
            oRed   <= 0;
            oGreen <= 0;
            oBlue  <= 0;
        end else begin
            if (!iVideo_On) begin
                // Text only (alarm mode)
                if (pixel_on2) begin
                    oRed   <= 0;
                    oGreen <= GREEN;
                    oBlue  <= 0;
                end else begin
                    oRed   <= BLACK;
                    oGreen <= BLACK;
                    oBlue  <= BLACK;
                end
            end else begin
                // Video + overlay
                if (pixel_on) begin
                    oRed   <= RED;
                    oGreen <= 0;
                    oBlue  <= 0;
						  
                end else if (video_region) begin
                    oRed   <= iRed;
                    oGreen <= iGreen;
                    oBlue  <= iBlue;
                end else begin
							oRed <= BLACK;
							oGreen <= BLACK;
							oBlue <= BLACK;
					 end
            end
        end
    end

endmodule
 
